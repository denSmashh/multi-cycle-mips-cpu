module cpu_top (
     input logic clk,
     input logic RSTn
     
);
    
    
    
endmodule
